`define NUM_OF_DUTS  1
`define NUM_OF_TRANS 4
